library verilog;
use verilog.vl_types.all;
entity sisc_tb is
    generic(
        tclk            : real    := 10.000000
    );
end sisc_tb;
